SHA512 (spice-0.15.1.tar.bz2) = 362ab2f0b483911830693834515e1d331a6b929c5c63fd4522e843c42bbb7d8a52510d60f5f17d175dd2617c9621630f6a81f3ff7dce11dc28e6fb135e60fa86
SHA512 (spice-0.15.1.tar.bz2.sig) = f53cd11edc73ca04a8518f412680c2afe27d2500e87284c17840d6ed0c8cb0d9ed71bc848b8bbaa04dda825ff93fa1f781ea496622a5440e5ccbeedde13cbc5c
SHA512 (victortoso-E37A484F.keyring) = 091755da8a358c8c8ebd3b5443b4b5eb3c260afed943454c085d48c973de6a42763547c321c64e4da5c1b2983ad0c5146aaeddeb1d54ef414f7e6a530a3bf14a
